----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/05/2024 10:30:24 PM
-- Design Name: 
-- Module Name: charLib - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity charLib is
    Port ( clka : in STD_LOGIC;
           addra : in STD_LOGIC_VECTOR (10 downto 0);
           douta : out STD_LOGIC_VECTOR (7 downto 0));
end charLib;

architecture Behavioral of charLib is

type ARR is Array (0 to 1023) of std_logic_vector (7 downto 0); 
signal characterlibrary :ARR := (
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
	x"00",x"00",x"00",x"5f",x"00",x"00",x"00",x"00",
	x"00",x"00",x"03",x"00",x"03",x"00",x"00",x"00",
	x"64",x"3c",x"26",x"64",x"3c",x"26",x"24",x"00",
	x"26",x"49",x"49",x"7f",x"49",x"49",x"32",x"00",
	x"42",x"25",x"12",x"08",x"24",x"52",x"21",x"00",
	x"20",x"50",x"4e",x"55",x"22",x"58",x"28",x"00",
	x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",
	x"00",x"00",x"1c",x"22",x"41",x"00",x"00",x"00",
	x"00",x"00",x"00",x"41",x"22",x"1c",x"00",x"00",
	x"00",x"15",x"15",x"0e",x"0e",x"15",x"15",x"00",
	x"00",x"08",x"08",x"3e",x"08",x"08",x"00",x"00",
	x"00",x"00",x"00",x"50",x"30",x"00",x"00",x"00",
	x"00", x"08", x"08", x"08", x"08", x"08", x"00", x"00",
    x"00", x"00", x"00", x"40", x"00", x"00", x"00", x"00",
x"40", x"20", x"10", x"08", x"04", x"02", x"01", x"00",
x"00", x"3E", x"41", x"41", x"41", x"3E", x"00", x"00",
x"00", x"00", x"41", x"7F", x"40", x"00", x"00", x"00",
x"00", x"42", x"61", x"51", x"49", x"6E", x"00", x"00",

	x"00", x"22", x"41", x"49", x"49", x"36", x"00", x"00",
x"00", x"18", x"14", x"12", x"7F", x"10", x"00", x"00",
x"00", x"27", x"49", x"49", x"49", x"71", x"00", x"00",
x"00", x"3C", x"4A", x"49", x"48", x"70", x"00", x"00",
x"00", x"43", x"21", x"11", x"0D", x"03", x"00", x"00",
x"00", x"36", x"49", x"49", x"49", x"36", x"00", x"00",
x"00", x"06", x"09", x"49", x"29", x"1E", x"00", x"00",
x"00", x"00", x"00", x"12", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"52", x"30", x"00", x"00", x"00",
x"00", x"00", x"08", x"14", x"14", x"22", x"00", x"00",
x"00", x"14", x"14", x"14", x"14", x"14", x"14", x"00",
x"00", x"00", x"22", x"14", x"14", x"08", x"00", x"00",
x"00", x"02", x"01", x"59", x"05", x"02", x"00", x"00",
x"3E", x"41", x"5D", x"55", x"4D", x"51", x"2E", x"00",
x"40", x"7C", x"4A", x"09", x"4A", x"7C", x"40", x"00",
x"41", x"7F", x"49", x"49", x"49", x"49", x"36", x"00",
x"1C", x"22", x"41", x"41", x"41", x"41", x"22", x"00",
x"41", x"7F", x"41", x"41", x"41", x"22", x"1C", x"00",
x"41", x"7F", x"49", x"49", x"5D", x"41", x"63", x"00",
x"41", x"7F", x"49", x"09", x"1D", x"01", x"03", x"00",
x"1C", x"22", x"41", x"49", x"49", x"3A", x"08", x"00",
x"41", x"7F", x"08", x"08", x"08", x"7F", x"41", x"00",
x"00", x"41", x"41", x"7F", x"41", x"41", x"00", x"00",
x"30", x"40", x"41", x"41", x"3F", x"01", x"01", x"00",
x"41", x"7F", x"08", x"0C", x"12", x"61", x"41", x"00",
x"41", x"7F", x"41", x"40", x"40", x"40", x"60", x"00",
x"41", x"7F", x"42", x"0C", x"42", x"7F", x"41", x"00",
x"41", x"7F", x"42", x"0C", x"11", x"7F", x"01", x"00",
x"1C", x"22", x"41", x"41", x"41", x"22", x"1C", x"00",
x"41", x"7F", x"49", x"09", x"09", x"09", x"06", x"00",
x"0C", x"12", x"21", x"21", x"61", x"52", x"4C", x"00",
x"41", x"7F", x"09", x"09", x"19", x"69", x"46", x"00",
x"66", x"49", x"49", x"49", x"49", x"49", x"33", x"00",
x"03", x"01", x"41", x"7F", x"41", x"01", x"03", x"00",
x"01", x"3F", x"41", x"40", x"41", x"3F", x"01", x"00",
x"01", x"0F", x"31", x"40", x"31", x"0F", x"01", x"00",
x"01", x"1F", x"61", x"14", x"61", x"1F", x"01", x"00",
x"41", x"41", x"36", x"08", x"36", x"41", x"41", x"00",
x"01", x"03", x"44", x"78", x"44", x"03", x"01", x"00",
x"43", x"61", x"51", x"49", x"45", x"43", x"61", x"00",
x"00", x"00", x"7F", x"41", x"41", x"00", x"00", x"00",
x"01", x"02", x"04", x"08", x"10", x"20", x"40", x"00",
x"00", x"00", x"41", x"41", x"7F", x"00", x"00", x"00",
x"00", x"04", x"02", x"01", x"01", x"02", x"04", x"00",
x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"00",
x"00", x"01", x"02", x"00", x"00", x"00", x"00", x"00",
x"00", x"34", x"4A", x"4A", x"4A", x"3C", x"40", x"00",
x"00", x"41", x"3F", x"48", x"48", x"48", x"30", x"00",
x"00", x"3C", x"42", x"42", x"42", x"24", x"00", x"00",
x"00", x"30", x"48", x"48", x"49", x"3F", x"40", x"00",
x"00", x"3C", x"4A", x"4A", x"4A", x"2C", x"00", x"00",
x"00", x"00", x"48", x"7E", x"49", x"09", x"00", x"00",
x"00", x"26", x"49", x"49", x"49", x"3F", x"01", x"00",
x"41", x"7F", x"48", x"04", x"44", x"78", x"40", x"00",
x"00", x"00", x"44", x"7D", x"40", x"00", x"00", x"00",
x"00", x"00", x"40", x"44", x"3D", x"00", x"00", x"00",
x"41", x"7F", x"10", x"18", x"24", x"42", x"42", x"00",
x"00", x"40", x"41", x"7F", x"40", x"40", x"00", x"00",
x"42", x"7E", x"02", x"7C", x"02", x"7E", x"40", x"00",
x"42", x"7E", x"44", x"02", x"42", x"7C", x"40", x"00",
x"00", x"3C", x"42", x"42", x"42", x"3C", x"00", x"00",
x"00", x"41", x"7F", x"49", x"09", x"09", x"06", x"00",
x"00", x"06", x"09", x"09", x"49", x"7F", x"41", x"00",
x"00", x"42", x"7E", x"44", x"02", x"02", x"04", x"00",
x"00", x"64", x"4A", x"4A", x"4A", x"36", x"00", x"00",
x"00", x"04", x"3F", x"44", x"44", x"20", x"00", x"00",
x"00", x"02", x"3E", x"40", x"40", x"22", x"7E", x"40",
x"02", x"0E", x"32", x"40", x"32", x"0E", x"02", x"00",
x"02", x"1E", x"62", x"18", x"62", x"1E", x"02", x"00",
x"42", x"62", x"14", x"08", x"14", x"62", x"42", x"00",
x"01", x"43", x"45", x"38", x"05", x"03", x"01", x"00",
x"00", x"46", x"62", x"52", x"4A", x"46", x"62", x"00",
x"00", x"00", x"08", x"36", x"41", x"00", x"00", x"00",
x"00", x"00", x"00", x"7F", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"41", x"36", x"08", x"00", x"00",
x"00", x"18", x"08", x"08", x"10", x"10", x"18", x"00",
x"AA", x"55", x"AA", x"55", x"AA", x"55", x"AA", x"55");


begin

process(clka)
begin 

    if(rising_edge(clka)) then 
        
        douta <= characterlibrary( to_integer(unsigned(addra))); 
        
    end if; 
    
end process;  

end Behavioral;
